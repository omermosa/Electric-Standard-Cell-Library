*** SPICE deck for cell Complex_1_sim{sch} from library Complex
*** Created on Mon Apr 13, 2020 23:27:55
*** Last revised on Sat Apr 18, 2020 17:31:25
*** Written on Sun Apr 19, 2020 04:01:57 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Complex__Complex_1 FROM CELL Complex_1{sch}
.SUBCKT Complex__Complex_1 f w x y z
** GLOBAL gnd
** GLOBAL vdd
** GLOBAL x
** GLOBAL y
** GLOBAL z
** GLOBAL w
Mnmos@0 net@5 y gnd gnd NMOS L=0.36U W=2.34U
Mnmos@1 f x net@5 gnd NMOS L=0.36U W=2.34U
Mnmos@2 net@4 z gnd gnd NMOS L=0.36U W=2.34U
Mnmos@4 f w net@4 gnd NMOS L=0.36U W=2.34U
Mpmos@0 net@20 x f vdd PMOS L=0.36U W=4.32U
Mpmos@1 net@20 y f vdd PMOS L=0.36U W=4.32U
Mpmos@2 vdd w net@20 vdd PMOS L=0.36U W=4.32U
Mpmos@3 vdd z net@20 vdd PMOS L=0.36U W=4.32U
.ENDS Complex__Complex_1

.global gnd vdd x y z w

*** TOP LEVEL CELL: Complex_1_sim{sch}
XComplex_@0 f vdd gnd gnd z Complex__Complex_1

* Spice Code nodes in cell cell 'Complex_1_sim{sch}'
vdd vdd 0 dc 3.3
vz z 0 DC pulse 0 3.3  1n .001n .001n 5n 10n
cload f 0 16fF
.tran 0 100n
.measure tdpr trig v(z) val=1.65 fall =1 TARG v(f) val=1.65 rise=1
.measure tdpf trig v(z) val=1.65 rise =1 TARG v(f) val=1.65 fall=1
.measure trise trig v(f) val=0.66 rise =1 TARG v(f) val=2.64 rise=1
.measure tfall trig v(f) val=2.64 fall =1 TARG v(f) val=0.66 fall=1
.include D:\AUC\Spring_20\DD2\Electric\scmos18.txt
.END
