*** SPICE deck for cell tristate_inv_1_sim{sch} from library Tristate_Inv
*** Created on Fri Apr 17, 2020 20:56:21
*** Last revised on Fri Apr 17, 2020 22:06:14
*** Written on Sun Apr 19, 2020 04:14:40 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Tristate_Inv__tristate_inv_1 FROM CELL tristate_inv_1{sch}
.SUBCKT Tristate_Inv__tristate_inv_1 En En_ In OUT
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 OUT En net@13 gnd NMOS L=0.36U W=1.8U
Mnmos@2 net@13 In gnd gnd NMOS L=0.36U W=1.8U
Mpmos@1 vdd In net@15 vdd PMOS L=0.36U W=5.04U
Mpmos@2 net@15 En_ OUT vdd PMOS L=0.36U W=5.04U
.ENDS Tristate_Inv__tristate_inv_1

.global gnd vdd

*** TOP LEVEL CELL: tristate_inv_1_sim{sch}
Xtristate@0 vdd gnd in out Tristate_Inv__tristate_inv_1

* Spice Code nodes in cell cell 'tristate_inv_1_sim{sch}'
vdd vdd 0 dc 3.3
vin in 0 DC pulse 0 3.3  1n .001n .001n 5n 10n
cload out 0 16fF
.tran 0 100n
.measure tdpr trig v(in) val=1.65 fall =1 TARG v(out) val=1.65 rise=1
.measure tdpf trig v(in) val=1.65 rise =1 TARG v(out) val=1.65 fall=1
.measure trise trig v(out) val=0.66 rise =1 TARG v(out) val=2.64 rise=1
.measure tfall trig v(out) val=2.64 fall =1 TARG v(out) val=0.66 fall=1
.include D:\AUC\Spring_20\DD2\Electric\scmos18.txt
.END
