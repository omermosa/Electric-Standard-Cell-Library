*** SPICE deck for cell sim_Inverter_1{sch} from library Inverter
*** Created on Fri Apr 17, 2020 04:37:34
*** Last revised on Fri Apr 17, 2020 05:01:37
*** Written on Fri Apr 17, 2020 05:06:39 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Inverter__Inverter_1 FROM CELL Inverter:Inverter_1{sch}
.SUBCKT Inverter__Inverter_1 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.36U W=0.9U
Mpmos@0 vdd in out vdd P L=0.36U W=2.16U
.ENDS Inverter__Inverter_1

.global gnd vdd

*** TOP LEVEL CELL: Inverter:sim_Inverter_1{sch}
XInverter@0 in out Inverter__Inverter_1

* Spice Code nodes in cell cell 'Inverter:sim_Inverter_1{sch}'
vdd vdd 0 dc 3.3
vin in 0 DC pulse 0 3.3  1n 1.333n 1.333n 5n 12.667n
cload out 0 128fF
.tran 0 100n
.measure tdpr trig v(in) val=1.65 fall =1 TARG v(out) val=1.65 rise=1
.measure tdpf trig v(in) val=1.65 rise =1 TARG v(out) val=1.65 fall=1
.measure trise trig v(out) val=0.66 rise =1 TARG v(out) val=2.64 rise=1
.measure tfall trig v(out) val=2.64 fall =1 TARG v(out) val=0.66 fall=1
.include scmos18.txt
.END
